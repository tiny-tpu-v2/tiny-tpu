module accumulator (
)

endmodule