module dump();
initial begin
    $dumpfile("float32_adder.vcd");
    $dumpvars(0, float32_adder);
end
endmodule