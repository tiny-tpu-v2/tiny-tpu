`timescale 1ns/1ps
`default_nettype none

module vector_unit (
    

);


endmodule